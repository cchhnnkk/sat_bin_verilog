
int nb = 3;
int cmax = 8;
int vmax = 8;

int cbin[24][8] = '{
	//bin 1
	'{1, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},

	//bin 2
	'{2, 0, 1, 0, 0, 0, 0, 0},
	'{0, 2, 0, 1, 0, 0, 0, 0},
	'{0, 0, 2, 0, 2, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},

	//bin 3
	'{1, 0, 2, 0, 2, 0, 0, 0},
	'{0, 2, 0, 1, 1, 0, 0, 0},
	'{0, 2, 0, 0, 2, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0}
};

int vbin[24] = '{
	//bin 1
	1, 0, 0, 0, 0, 0, 0, 0,
	//bin 2
	2, 3, 4, 5, 6, 0, 0, 0,
	//bin 3
	1, 2, 5, 6, 7, 0, 0, 0
};


