module sat_engine #(
	parameter ACTIVITY_BASE_ADDR = 0,
	parameter MEM_DATA_WIDTH = 512,
	parameter VAR_WIDTH = 15,
	parameter VALUE_ADDR_WIDTH = VAR_WIDTH,
	parameter LEVEL_DATA_WIDTH = 9,
	parameter LEVEL_ADDR_WIDTH = VAR_WIDTH,
	parameter ACTIVITY_DATA_WIDTH = 16,
	parameter ACTIVITY_ADDR_WIDTH = VAR_WIDTH,
 )(
	wire clk,
	wire rst,
);




endmodule
