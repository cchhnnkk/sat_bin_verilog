
int nb1 = 3;
int cmax1 = 8;
int vmax1 = 8;

int cbin1[24][8] = '{
	//bin 1
	'{1, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},

	//bin 2
	'{2, 0, 1, 0, 0, 0, 0, 0},
	'{0, 2, 0, 1, 0, 0, 0, 0},
	'{0, 0, 2, 0, 2, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},

	//bin 3
	'{1, 0, 2, 0, 2, 0, 0, 0},
	'{0, 2, 0, 1, 1, 0, 0, 0},
	'{0, 2, 0, 0, 2, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0},
	'{0, 0, 0, 0, 0, 0, 0, 0}
};

int vbin1[24] = '{
	//bin 1
	1, 0, 0, 0, 0, 0, 0, 0,
	//bin 2
	2, 3, 4, 5, 6, 0, 0, 0,
	//bin 3
	1, 2, 5, 6, 7, 0, 0, 0
};

task bm_test_case1();
    nb = nb1;
    cmax = cmax1;
    vmax = vmax1;
    cbin = cbin1;
    vbin = vbin1;
    run_test_case();
endtask

